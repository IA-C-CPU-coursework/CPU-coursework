

module mips_decoder_tb()