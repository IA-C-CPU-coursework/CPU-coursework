module mips_cpu_alu_control(
input ALUOp,
input FuncCode,
output ALUControl
);

